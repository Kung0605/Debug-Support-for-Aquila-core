module cdc_4phase #(
  parameter type T = logic,
  parameter bit DECOUPLED = 1'b1,
  parameter bit SEND_RESET_MSG = 1'b0,
  parameter T RESET_MSG = T'('0)
)(
  input  logic src_rst_ni,
  input  logic src_clk_i,
  input  T     src_data_i,
  input  logic src_valid_i,
  output logic src_ready_o,

  input  logic dst_rst_ni,
  input  logic dst_clk_i,
  output T     dst_data_o,
  output logic dst_valid_o,
  input  logic dst_ready_i
);

  // Asynchronous handshake signals.
  (* dont_touch = "true" *) logic async_req;
  (* dont_touch = "true" *) logic async_ack;
  (* dont_touch = "true" *) T async_data;

  // The sender in the source domain.
  cdc_4phase_src #(
    .T(T),
    .DECOUPLED(DECOUPLED),
    .SEND_RESET_MSG(SEND_RESET_MSG),
    .RESET_MSG(RESET_MSG)
  ) i_src (
    .rst_ni       ( src_rst_ni  ),
    .clk_i        ( src_clk_i   ),
    .data_i       ( src_data_i  ),
    .valid_i      ( src_valid_i ),
    .ready_o      ( src_ready_o ),
    .async_req_o  ( async_req   ),
    .async_ack_i  ( async_ack   ),
    .async_data_o ( async_data  )
  );

  // The receiver in the destination domain.
  cdc_4phase_dst #(.T(T), .DECOUPLED(DECOUPLED)) i_dst (
    .rst_ni       ( dst_rst_ni  ),
    .clk_i        ( dst_clk_i   ),
    .data_o       ( dst_data_o  ),
    .valid_o      ( dst_valid_o ),
    .ready_i      ( dst_ready_i ),
    .async_req_i  ( async_req   ),
    .async_ack_o  ( async_ack   ),
    .async_data_i ( async_data  )
  );
endmodule


/// Half of the 4-phase clock domain crossing located in the source domain.
module cdc_4phase_src #(
  parameter type T = logic,
  parameter int unsigned SYNC_STAGES = 2,
  parameter bit DECOUPLED = 1'b1,
  parameter bit SEND_RESET_MSG = 1'b0,
  parameter T RESET_MSG = T'('0)
)(
  input  logic rst_ni,
  input  logic clk_i,
  input  T     data_i,
  input  logic valid_i,
  output logic ready_o,
  output logic async_req_o,
  input  logic async_ack_i,
  output T     async_data_o
);

  (* dont_touch = "true" *)
  logic  req_src_d, req_src_q;
  (* dont_touch = "true" *)
  T data_src_d, data_src_q;
  (* dont_touch = "true" *)
  logic  ack_synced;

  typedef enum logic[1:0] {S_IDLE, S_WAIT_ACK_ASSERT, S_WAIT_ACK_DEASSERT} state_e;
  state_e src_state_d, src_state_q;

  // Synchronize the async ACK
  reg  [SYNC_STAGES-1:0] ack_synced_reg;

  always_ff @(posedge clk_i, negedge rst_ni) begin 
    if (~rst_ni)
      ack_synced_reg <= 0;
    else 
      ack_synced_reg <= {ack_synced_reg[SYNC_STAGES-2:0], async_ack_i};
  end

  assign ack_synced = ack_synced_reg[SYNC_STAGES-1];


  // FSM for the 4-phase handshake
  always_comb begin
    src_state_d    = src_state_q;
    req_src_d  = 1'b0;
    data_src_d = data_src_q;
    ready_o    = 1'b0;
    case (src_state_q)
      S_IDLE: begin
        // If decoupling is disabled, defer assertion of ready until the
        // handshake with the dst is completed
        if (DECOUPLED) begin
          ready_o = 1'b1;
        end else begin
          ready_o = 1'b0;
        end
        // Sample a new item when the valid signal is asserted.
        if (valid_i) begin
          data_src_d = data_i;
          req_src_d  = 1'b1;
          src_state_d = S_WAIT_ACK_ASSERT;
        end
      end
      S_WAIT_ACK_ASSERT: begin
        req_src_d = 1'b1;
        if (ack_synced == 1'b1) begin
          req_src_d = 1'b0;
          src_state_d   = S_WAIT_ACK_DEASSERT;
        end
      end
      S_WAIT_ACK_DEASSERT: begin
        if (ack_synced == 1'b0) begin
          src_state_d = S_IDLE;
          if (!DECOUPLED) begin
            ready_o = 1'b1;
          end
        end
      end
      default: begin
        src_state_d = S_IDLE;
      end
    endcase
  end

  always_ff @(posedge clk_i, negedge rst_ni) begin
    if (!rst_ni) begin
      src_state_q <= S_IDLE;
    end else begin
      src_state_q <= src_state_d;
    end
  end

  // Sample the data and the request signal to filter combinational glitches
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      if (SEND_RESET_MSG) begin
        req_src_q  <= 1'b1;
        data_src_q <= RESET_MSG;
      end else begin
        req_src_q  <= 1'b0;
        data_src_q <= T'('0);
      end
    end else begin
      req_src_q  <= req_src_d;
      data_src_q <= data_src_d;
    end
  end

  // Async output assignments.
  assign async_req_o = req_src_q;
  assign async_data_o = data_src_q;

endmodule


/// Half of the 4-phase clock domain crossing located in the destination domain.
module cdc_4phase_dst #(
  parameter type T = logic,
  parameter int unsigned SYNC_STAGES = 2,
  parameter bit DECOUPLED = 1
)(
  input  logic rst_ni,
  input  logic clk_i,
  output T     data_o,
  output logic valid_o,
  input  logic ready_i,
  input  logic async_req_i,
  output logic async_ack_o,
  input  T     async_data_i
);

  (* dont_touch = "true" *)
  logic  ack_dst_d, ack_dst_q;
  (* dont_touch = "true" *)
  logic  req_synced;

  logic  data_valid;

  logic  output_ready;


  typedef enum logic[1:0] {D_IDLE, D_WAIT_DOWNSTREAM_ACK, D_WAIT_REQ_DEASSERT} state_e;
  state_e dst_state_d, dst_state_q;
  
  //Synchronize the request
  reg  [SYNC_STAGES-1:0] req_synced_reg;

  always_ff @(posedge clk_i, negedge rst_ni) begin 
    if (~rst_ni)
      req_synced_reg <= 0;
    else 
      req_synced_reg <= {req_synced_reg[SYNC_STAGES-2:0], async_req_i};
  end

  assign req_synced = req_synced_reg[SYNC_STAGES-1];


  // FSM for the 4-phase handshake
  always_comb begin
    dst_state_d    = dst_state_q;
    data_valid = 1'b0;
    ack_dst_d  = 1'b0;

    case (dst_state_q)
      D_IDLE: begin
        // Sample the data upon a new request and transition to the next state
        if (req_synced == 1'b1) begin
          data_valid = 1'b1;
          if (output_ready == 1'b1) begin
            dst_state_d = D_WAIT_REQ_DEASSERT;
          end else begin
            dst_state_d = D_WAIT_DOWNSTREAM_ACK;
          end
        end
      end

      D_WAIT_DOWNSTREAM_ACK: begin
        data_valid       = 1'b1;
        if (output_ready == 1'b1) begin
          dst_state_d    = D_WAIT_REQ_DEASSERT;
          ack_dst_d  = 1'b1;
        end
      end

      D_WAIT_REQ_DEASSERT: begin
        ack_dst_d = 1'b1;
        if (req_synced == 1'b0) begin
          ack_dst_d = 1'b0;
          dst_state_d   = D_IDLE;
        end
      end

      default: begin
        dst_state_d = D_IDLE;
      end
    endcase
  end

  always_ff @(posedge clk_i, negedge rst_ni) begin
    if (!rst_ni) begin
      dst_state_q <= D_IDLE;
    end else begin
      dst_state_q <= dst_state_d;
    end
  end

  // Filter glitches on ack signal before sending it through the asynchronous channel
  always_ff @(posedge clk_i, negedge rst_ni) begin
    if (!rst_ni) begin
      ack_dst_q <= 1'b0;
    end else begin
      ack_dst_q <= ack_dst_d;
    end
  end

  assign valid_o      = data_valid;
  assign output_ready = ready_i;
  assign data_o       = async_data_i;

  // Output assignments.
  assign async_ack_o = ack_dst_q;

endmodule